module INSTMEM(PC,inst,clk);
	input[31:0] PC;
	input clk;
	output[31:0] inst;
	reg[31:0] inst;
	reg[31:0] memory[0:31];
	integer mem;
	initial begin
    	memory[0] = 32'b00000000000000000000000000000000;  
    	memory[1] = 32'b00000000000000000000000000000000;  
    	memory[2] = 32'b00000000000000000000000000000000;  
    	memory[3] = 32'b10001100000100010000000000001000;  // lw  $s1($17), 8($0)
    	memory[4] = 32'b10001100000100100000000000000100;  // lw  $s2($18), 4($0)
    	memory[5] = 32'b00000010001100100100000000100000;  // add $t0($8), $s1($17), $s2($18)
    	memory[6] = 32'b00000000000000000000000000000000;  // nop
    	memory[7] = 32'b00000000000000000000000000000000;  // nop
    	memory[8] = 32'b00000000000000000000000000000000;  // nop
    	memory[9] = 32'b00000000000000000000000000000000;  // nop
    	memory[10]= 32'b00000000000000000000000000000000;  // nop
    	memory[11]= 32'b00000000000000000000000000000000;  // nop
    	memory[12]= 32'b00000000000000000000000000000000;  // nop
    	memory[13]= 32'b00000000000000000000000000000000;  // nop
    	memory[14]= 32'b00000000000000000000000000000000;  // nop
    	memory[15]= 32'b00000000000000000000000000000000;  // nop
    	memory[16]= 32'b00000000000000000000000000000000;  // nop
    	memory[17]= 32'b00000000000000000000000000000000;  // nop
    	memory[18]= 32'b00000000000000000000000000000000;  // nop 
    	memory[19]= 32'b00000000000000000000000000000000;  // nop
    	memory[20]= 32'b00000000000000000000000000000000;  // nop
    	memory[21]= 32'b00000000000000000000000000000000;  // nop
    	memory[22]= 32'b00000000000000000000000000000000;  // nop
    	memory[23]= 32'b00000000000000000000000000000000;  // nop
    	memory[24]= 32'b00000000000000000000000000000000;  // nop
    	memory[25]= 32'b00000000000000000000000000000000;  // nop
    	memory[26]= 32'b00000000000000000000000000000000;  // nop
    	memory[27]= 32'b00000000000000000000000000000000;  // nop
    	memory[28]= 32'b00000000000000000000000000000000;  // nop 
    	memory[29]= 32'b00000000000000000000000000000000;  // nop
    	memory[30]= 32'b00000000000000000000000000000000;  // nop
    	memory[31]= 32'b00000000000000000000000000000000;
	end
	always@(posedge clk)
	begin
	mem = PC[31:0];
	inst = memory[mem];
	end
endmodule

/*module testINST;
	reg clk,reset;
	reg[31:0] PC;
	wire[31:0] out;
	wire[31:0] out1;
	PC pc(out,clk,reset);
	INSTMEM I(out,out1,clk);
	initial
	begin
		$monitor($time,"PCout=%b inst=%b",out,out1);
		#0 reset = 1'b1;clk=1'b0;
		#10 reset = 1'b0;
	end
	initial
	begin
	repeat(1000)
	#1 clk = ~clk;
	end
endmodule*/
