module SCDdatapath(ALUout,PC,reset,clk);
	input clk,reset;
	input[31:0] PC;
	output[31:0] aluout;
endmodule;
	
	
	
	
	
	
	
	
	
	
	
	
