module full_adder();
endmodule

module item();
endmodule
